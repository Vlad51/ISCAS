
module c432 ( N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, 
        N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, 
        N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, 
        N421, N430, N431, N432 );
  input N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47,
         N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92,
         N95, N99, N102, N105, N108, N112, N115;
  output N223, N329, N370, N421, N430, N431, N432;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318;

  NAND2_X2 U98 ( .A1(n120), .A2(n121), .ZN(n97) );
  AND2_X2 U99 ( .A1(n97), .A2(n98), .ZN(n286) );
  AND2_X2 U100 ( .A1(n99), .A2(n262), .ZN(n98) );
  INV_X1 U101 ( .A(N40), .ZN(n99) );
  NOR2_X2 U102 ( .A1(n305), .A2(n304), .ZN(n311) );
  INV_X4 U103 ( .A(n271), .ZN(n237) );
  INV_X4 U104 ( .A(n303), .ZN(n299) );
  NOR2_X2 U105 ( .A1(n288), .A2(N66), .ZN(n289) );
  INV_X8 U106 ( .A(n298), .ZN(n120) );
  OAI22_X4 U107 ( .A1(n139), .A2(N102), .B1(n138), .B2(N89), .ZN(n144) );
  INV_X4 U108 ( .A(N108), .ZN(n139) );
  INV_X1 U109 ( .A(n161), .ZN(n100) );
  INV_X4 U110 ( .A(n294), .ZN(n161) );
  INV_X1 U111 ( .A(n314), .ZN(n317) );
  AND2_X2 U112 ( .A1(n101), .A2(n262), .ZN(n170) );
  NOR2_X1 U113 ( .A1(N40), .A2(n168), .ZN(n101) );
  NAND2_X4 U114 ( .A1(n164), .A2(N30), .ZN(n165) );
  NAND2_X2 U115 ( .A1(n112), .A2(n179), .ZN(n180) );
  NAND2_X2 U116 ( .A1(n210), .A2(N17), .ZN(n211) );
  INV_X4 U117 ( .A(n211), .ZN(n251) );
  NOR2_X4 U118 ( .A1(n307), .A2(N115), .ZN(n308) );
  OAI21_X4 U119 ( .B1(n116), .B2(n297), .A(n103), .ZN(n307) );
  INV_X1 U120 ( .A(n127), .ZN(n102) );
  INV_X2 U121 ( .A(n102), .ZN(n103) );
  NOR2_X1 U122 ( .A1(n180), .A2(n189), .ZN(n117) );
  NAND2_X4 U123 ( .A1(n265), .A2(n262), .ZN(n169) );
  INV_X8 U124 ( .A(n165), .ZN(n262) );
  OAI22_X4 U125 ( .A1(n161), .A2(n193), .B1(n160), .B2(n208), .ZN(n104) );
  NAND2_X4 U126 ( .A1(n150), .A2(N37), .ZN(n177) );
  INV_X8 U127 ( .A(n105), .ZN(n110) );
  NOR2_X2 U128 ( .A1(n287), .A2(N53), .ZN(n290) );
  BUF_X16 U129 ( .A(n138), .Z(n105) );
  INV_X2 U130 ( .A(n276), .ZN(n106) );
  INV_X2 U131 ( .A(n106), .ZN(n107) );
  INV_X8 U132 ( .A(n250), .ZN(n257) );
  INV_X1 U133 ( .A(n116), .ZN(n108) );
  INV_X2 U134 ( .A(n283), .ZN(n264) );
  INV_X2 U135 ( .A(n206), .ZN(n160) );
  INV_X4 U136 ( .A(n274), .ZN(n247) );
  NOR2_X2 U137 ( .A1(n267), .A2(n276), .ZN(n268) );
  INV_X4 U138 ( .A(N430), .ZN(n316) );
  AOI21_X2 U139 ( .B1(n270), .B2(n269), .A(n268), .ZN(N432) );
  INV_X8 U140 ( .A(n180), .ZN(n240) );
  NOR2_X1 U141 ( .A1(n220), .A2(n213), .ZN(n218) );
  NAND2_X2 U142 ( .A1(n126), .A2(n182), .ZN(n183) );
  NOR2_X4 U143 ( .A1(n104), .A2(n184), .ZN(n185) );
  BUF_X16 U144 ( .A(n251), .Z(n125) );
  NAND2_X4 U145 ( .A1(n128), .A2(n167), .ZN(n172) );
  NAND2_X4 U146 ( .A1(n242), .A2(n240), .ZN(n190) );
  OAI22_X4 U147 ( .A1(n163), .A2(n213), .B1(n162), .B2(n216), .ZN(n184) );
  OAI22_X4 U148 ( .A1(n223), .A2(n209), .B1(n222), .B2(n208), .ZN(n219) );
  NAND2_X4 U149 ( .A1(n231), .A2(n229), .ZN(n222) );
  BUF_X16 U150 ( .A(n232), .Z(n109) );
  INV_X4 U151 ( .A(n215), .ZN(n232) );
  NAND2_X2 U152 ( .A1(n250), .A2(N27), .ZN(n260) );
  NOR2_X4 U153 ( .A1(n249), .A2(n248), .ZN(n270) );
  OAI22_X4 U154 ( .A1(n163), .A2(n213), .B1(n162), .B2(n216), .ZN(n111) );
  INV_X1 U155 ( .A(n155), .ZN(n112) );
  NAND2_X4 U156 ( .A1(n129), .A2(n128), .ZN(n113) );
  NAND2_X4 U157 ( .A1(n251), .A2(n212), .ZN(n220) );
  NAND2_X4 U158 ( .A1(n256), .A2(n254), .ZN(n198) );
  NAND2_X4 U159 ( .A1(n232), .A2(n235), .ZN(n221) );
  NAND4_X4 U160 ( .A1(n198), .A2(n190), .A3(n194), .A4(n192), .ZN(n186) );
  NOR2_X2 U161 ( .A1(n302), .A2(N79), .ZN(n305) );
  OAI21_X4 U162 ( .B1(n116), .B2(n244), .A(n243), .ZN(n302) );
  NAND2_X4 U163 ( .A1(n122), .A2(n262), .ZN(n283) );
  NAND2_X4 U164 ( .A1(n120), .A2(n121), .ZN(n122) );
  NAND2_X4 U165 ( .A1(n119), .A2(n238), .ZN(N370) );
  INV_X1 U166 ( .A(n267), .ZN(n114) );
  INV_X8 U167 ( .A(n188), .ZN(n115) );
  BUF_X16 U168 ( .A(n141), .Z(n124) );
  INV_X8 U169 ( .A(n318), .ZN(n266) );
  INV_X8 U170 ( .A(N370), .ZN(n246) );
  NAND2_X2 U171 ( .A1(n260), .A2(n261), .ZN(n277) );
  OAI21_X4 U172 ( .B1(n266), .B2(n235), .A(n234), .ZN(n236) );
  NOR2_X4 U173 ( .A1(n308), .A2(n309), .ZN(n310) );
  NOR3_X4 U174 ( .A1(n301), .A2(n300), .A3(n299), .ZN(n312) );
  OAI21_X4 U175 ( .B1(n298), .B2(n233), .A(n109), .ZN(n306) );
  NAND2_X4 U176 ( .A1(n226), .A2(n225), .ZN(n227) );
  NOR2_X1 U177 ( .A1(n221), .A2(n216), .ZN(n217) );
  INV_X8 U178 ( .A(n227), .ZN(n238) );
  NAND2_X2 U179 ( .A1(n242), .A2(n117), .ZN(n123) );
  INV_X8 U180 ( .A(n113), .ZN(n116) );
  NAND3_X2 U181 ( .A1(n123), .A2(n201), .A3(n200), .ZN(n118) );
  NOR3_X4 U182 ( .A1(n203), .A2(n115), .A3(n202), .ZN(n119) );
  OAI21_X4 U183 ( .B1(n172), .B2(n173), .A(n171), .ZN(n203) );
  NAND3_X2 U184 ( .A1(n149), .A2(n148), .A3(n147), .ZN(n150) );
  INV_X1 U185 ( .A(n263), .ZN(n121) );
  NAND2_X2 U186 ( .A1(N223), .A2(N89), .ZN(n214) );
  INV_X8 U187 ( .A(n183), .ZN(n243) );
  INV_X4 U188 ( .A(n124), .ZN(n130) );
  NOR2_X1 U189 ( .A1(n155), .A2(N60), .ZN(n156) );
  BUF_X4 U190 ( .A(N69), .Z(n126) );
  NAND2_X2 U191 ( .A1(n283), .A2(n284), .ZN(n282) );
  NAND3_X2 U192 ( .A1(n123), .A2(n201), .A3(n200), .ZN(n202) );
  NOR3_X2 U193 ( .A1(n219), .A2(n217), .A3(n218), .ZN(n226) );
  NOR2_X2 U194 ( .A1(n169), .A2(n175), .ZN(n166) );
  INV_X4 U195 ( .A(n277), .ZN(n267) );
  NOR2_X2 U196 ( .A1(n290), .A2(n289), .ZN(n291) );
  NOR2_X2 U197 ( .A1(n286), .A2(n285), .ZN(n292) );
  NOR3_X2 U198 ( .A1(n282), .A2(n281), .A3(n280), .ZN(n293) );
  NOR2_X2 U199 ( .A1(n194), .A2(n193), .ZN(n195) );
  INV_X4 U200 ( .A(n199), .ZN(n200) );
  NOR2_X2 U201 ( .A1(n198), .A2(n197), .ZN(n199) );
  NOR2_X2 U202 ( .A1(n306), .A2(N105), .ZN(n309) );
  INV_X4 U203 ( .A(N56), .ZN(n155) );
  INV_X4 U204 ( .A(N69), .ZN(n140) );
  NAND2_X2 U205 ( .A1(n205), .A2(n127), .ZN(n223) );
  NOR2_X2 U206 ( .A1(n259), .A2(n258), .ZN(n269) );
  NAND2_X4 U207 ( .A1(n230), .A2(n130), .ZN(n208) );
  INV_X1 U208 ( .A(n191), .ZN(n176) );
  NOR2_X2 U209 ( .A1(n253), .A2(n284), .ZN(n259) );
  INV_X8 U210 ( .A(n146), .ZN(n147) );
  OAI22_X4 U211 ( .A1(N37), .A2(n145), .B1(n155), .B2(N50), .ZN(n146) );
  NOR2_X2 U212 ( .A1(n139), .A2(n152), .ZN(n127) );
  INV_X2 U213 ( .A(n154), .ZN(n167) );
  NAND2_X2 U214 ( .A1(n156), .A2(n179), .ZN(n189) );
  NOR2_X2 U215 ( .A1(n192), .A2(n191), .ZN(n196) );
  NOR2_X4 U216 ( .A1(n104), .A2(n111), .ZN(n128) );
  INV_X2 U217 ( .A(n210), .ZN(n163) );
  NOR2_X4 U218 ( .A1(n154), .A2(n175), .ZN(n129) );
  NAND2_X2 U219 ( .A1(n271), .A2(n272), .ZN(n273) );
  INV_X2 U220 ( .A(n260), .ZN(n253) );
  NAND2_X4 U221 ( .A1(n153), .A2(n191), .ZN(n154) );
  NAND2_X2 U222 ( .A1(n110), .A2(n214), .ZN(n215) );
  NAND3_X4 U223 ( .A1(n187), .A2(n185), .A3(n186), .ZN(n188) );
  NAND2_X1 U224 ( .A1(n275), .A2(n274), .ZN(n278) );
  OAI21_X2 U225 ( .B1(n317), .B2(n316), .A(n315), .ZN(N421) );
  NAND2_X4 U226 ( .A1(n189), .A2(n158), .ZN(n175) );
  NOR3_X2 U227 ( .A1(n176), .A2(n175), .A3(n174), .ZN(n187) );
  NAND2_X1 U228 ( .A1(N8), .A2(n108), .ZN(n295) );
  NAND2_X4 U229 ( .A1(N223), .A2(N63), .ZN(n182) );
  NAND3_X2 U230 ( .A1(n126), .A2(n244), .A3(n182), .ZN(n191) );
  NAND2_X4 U231 ( .A1(n245), .A2(n243), .ZN(n192) );
  NOR2_X2 U232 ( .A1(n303), .A2(N92), .ZN(n304) );
  INV_X8 U233 ( .A(N82), .ZN(n141) );
  OAI211_X2 U234 ( .C1(n279), .C2(n278), .A(n114), .B(n107), .ZN(N431) );
  NAND2_X4 U235 ( .A1(n239), .A2(n238), .ZN(n250) );
  NAND2_X4 U236 ( .A1(n119), .A2(n238), .ZN(n318) );
  NAND2_X4 U237 ( .A1(n129), .A2(n128), .ZN(N329) );
  INV_X8 U238 ( .A(N329), .ZN(n298) );
  OAI22_X4 U239 ( .A1(n152), .A2(n209), .B1(n151), .B2(n197), .ZN(n174) );
  INV_X4 U240 ( .A(N11), .ZN(n131) );
  NAND2_X2 U241 ( .A1(N17), .A2(n131), .ZN(n136) );
  INV_X4 U242 ( .A(N1), .ZN(n132) );
  NAND2_X2 U243 ( .A1(N4), .A2(n132), .ZN(n135) );
  INV_X4 U244 ( .A(N24), .ZN(n133) );
  NAND2_X2 U245 ( .A1(N30), .A2(n133), .ZN(n134) );
  NAND3_X2 U246 ( .A1(n136), .A2(n135), .A3(n134), .ZN(n137) );
  INV_X4 U247 ( .A(n137), .ZN(n149) );
  INV_X4 U248 ( .A(N95), .ZN(n138) );
  NOR2_X4 U249 ( .A1(N63), .A2(n140), .ZN(n143) );
  NOR2_X4 U250 ( .A1(n141), .A2(N76), .ZN(n142) );
  NOR3_X4 U251 ( .A1(n144), .A2(n143), .A3(n142), .ZN(n148) );
  INV_X4 U252 ( .A(N43), .ZN(n145) );
  NAND3_X4 U253 ( .A1(n148), .A2(n149), .A3(n147), .ZN(N223) );
  NAND2_X2 U254 ( .A1(N102), .A2(n150), .ZN(n204) );
  INV_X4 U255 ( .A(n204), .ZN(n152) );
  INV_X4 U256 ( .A(N112), .ZN(n297) );
  NAND2_X2 U257 ( .A1(n297), .A2(N108), .ZN(n209) );
  INV_X4 U258 ( .A(n177), .ZN(n151) );
  INV_X4 U259 ( .A(N47), .ZN(n255) );
  NAND2_X2 U260 ( .A1(n255), .A2(N43), .ZN(n197) );
  INV_X4 U261 ( .A(n174), .ZN(n153) );
  NAND2_X2 U262 ( .A1(N223), .A2(N50), .ZN(n179) );
  INV_X4 U263 ( .A(N34), .ZN(n263) );
  NAND2_X2 U264 ( .A1(n263), .A2(N30), .ZN(n168) );
  INV_X4 U265 ( .A(n168), .ZN(n157) );
  NAND2_X2 U266 ( .A1(N24), .A2(N223), .ZN(n164) );
  NAND2_X2 U267 ( .A1(n157), .A2(n164), .ZN(n158) );
  NAND2_X2 U268 ( .A1(N1), .A2(N223), .ZN(n294) );
  INV_X4 U269 ( .A(N8), .ZN(n159) );
  NAND2_X2 U270 ( .A1(n159), .A2(N4), .ZN(n193) );
  NAND2_X2 U271 ( .A1(N223), .A2(N76), .ZN(n206) );
  INV_X4 U272 ( .A(N86), .ZN(n230) );
  NAND2_X2 U273 ( .A1(N223), .A2(N11), .ZN(n210) );
  INV_X4 U274 ( .A(N21), .ZN(n252) );
  NAND2_X2 U275 ( .A1(n252), .A2(N17), .ZN(n213) );
  INV_X4 U276 ( .A(n214), .ZN(n162) );
  INV_X4 U277 ( .A(N99), .ZN(n233) );
  NAND2_X2 U278 ( .A1(n233), .A2(n110), .ZN(n216) );
  INV_X4 U279 ( .A(N40), .ZN(n265) );
  INV_X4 U280 ( .A(n166), .ZN(n173) );
  INV_X4 U281 ( .A(n170), .ZN(n171) );
  INV_X4 U282 ( .A(N53), .ZN(n256) );
  NAND2_X2 U283 ( .A1(N43), .A2(n177), .ZN(n178) );
  INV_X4 U284 ( .A(n178), .ZN(n254) );
  INV_X4 U285 ( .A(N66), .ZN(n242) );
  INV_X4 U286 ( .A(N14), .ZN(n181) );
  NAND3_X2 U287 ( .A1(n294), .A2(N4), .A3(n181), .ZN(n194) );
  INV_X4 U288 ( .A(N79), .ZN(n245) );
  NOR2_X4 U289 ( .A1(n196), .A2(n195), .ZN(n201) );
  NOR3_X4 U290 ( .A1(n203), .A2(n115), .A3(n118), .ZN(n239) );
  INV_X4 U291 ( .A(N115), .ZN(n205) );
  INV_X4 U292 ( .A(N92), .ZN(n231) );
  NAND2_X2 U293 ( .A1(n130), .A2(n206), .ZN(n207) );
  INV_X4 U294 ( .A(n207), .ZN(n229) );
  INV_X4 U295 ( .A(N27), .ZN(n212) );
  INV_X4 U296 ( .A(N105), .ZN(n235) );
  NAND4_X2 U297 ( .A1(n223), .A2(n222), .A3(n221), .A4(n220), .ZN(n224) );
  NAND3_X2 U298 ( .A1(n129), .A2(n185), .A3(n224), .ZN(n225) );
  OAI21_X4 U299 ( .B1(n298), .B2(n230), .A(n229), .ZN(n303) );
  OAI21_X4 U300 ( .B1(n257), .B2(n231), .A(n299), .ZN(n271) );
  INV_X4 U301 ( .A(n306), .ZN(n234) );
  NOR2_X4 U302 ( .A1(n237), .A2(n236), .ZN(n249) );
  INV_X4 U303 ( .A(N60), .ZN(n241) );
  OAI21_X4 U304 ( .B1(n116), .B2(n241), .A(n240), .ZN(n288) );
  INV_X4 U305 ( .A(n288), .ZN(n281) );
  OAI21_X4 U306 ( .B1(n246), .B2(n242), .A(n281), .ZN(n274) );
  INV_X4 U307 ( .A(N73), .ZN(n244) );
  INV_X4 U308 ( .A(n302), .ZN(n300) );
  OAI21_X4 U309 ( .B1(n245), .B2(n246), .A(n300), .ZN(n272) );
  NOR2_X4 U310 ( .A1(n247), .A2(n272), .ZN(n248) );
  OAI21_X4 U311 ( .B1(n116), .B2(n252), .A(n125), .ZN(n284) );
  OAI21_X4 U312 ( .B1(n116), .B2(n255), .A(n254), .ZN(n287) );
  INV_X4 U313 ( .A(n287), .ZN(n280) );
  OAI21_X4 U314 ( .B1(n257), .B2(n256), .A(n280), .ZN(n275) );
  INV_X4 U315 ( .A(n275), .ZN(n258) );
  INV_X4 U316 ( .A(n284), .ZN(n261) );
  OAI21_X4 U317 ( .B1(n266), .B2(n265), .A(n264), .ZN(n276) );
  INV_X4 U318 ( .A(n273), .ZN(n279) );
  NOR2_X4 U319 ( .A1(n284), .A2(N27), .ZN(n285) );
  OAI211_X2 U320 ( .C1(n293), .C2(n318), .A(n292), .B(n291), .ZN(N430) );
  NAND2_X2 U321 ( .A1(N14), .A2(n318), .ZN(n296) );
  NAND4_X2 U322 ( .A1(n296), .A2(n295), .A3(N4), .A4(n100), .ZN(n314) );
  NAND2_X2 U323 ( .A1(n306), .A2(n307), .ZN(n301) );
  OAI211_X2 U324 ( .C1(n318), .C2(n312), .A(n311), .B(n310), .ZN(n313) );
  NAND2_X2 U325 ( .A1(n313), .A2(n314), .ZN(n315) );
endmodule

