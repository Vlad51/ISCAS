//Verilog
//testbench ISCAS-85 c432

`timescale 1 ns/ 1 ps //����������� ��������� ������������� (1 �����������) � ������������ ������������ (1 �����������) - ����� 1000 �������������

module test_c432_1(); //������ testbench ������

//���������� ��������������� ������� ��������
reg  tN1,tN4,tN8,tN11,tN14,tN17,tN21,tN24,tN27,tN30,
     tN34,tN37,tN40,tN43,tN47,tN50,tN53,tN56,tN60,tN63,
     tN66,tN69,tN73,tN76,tN79,tN82,tN86,tN89,tN92,tN95,
     tN99,tN102,tN105,tN108,tN112,tN115;

//���������� ��������������� �������� ��������
wire tN223,tN329,tN370,tN421,tN430,tN431,tN432;

//�������� ���������� testbench ������
c432 ts(tN1,tN4,tN8,tN11,tN14,tN17,tN21,tN24,tN27,tN30,
        tN34,tN37,tN40,tN43,tN47,tN50,tN53,tN56,tN60,tN63,
        tN66,tN69,tN73,tN76,tN79,tN82,tN86,tN89,tN92,tN95,
        tN99,tN102,tN105,tN108,tN112,tN115,
        tN223,tN329,tN370,tN421,tN430,tN431,tN432); 

//������������� ������������ ��������� � ������ test
initial begin: test

//��� ������ ������������ ��������� ����������

//��������� ������ ���������� ������������� (scientific data)
$display("���������� ������������� ISCAS-85 c432:");

//����������� ������� ������� �������������
$timeformat(-9,1,"ns",8);

//����������� ������ ������� ������ � ���������� � ������� �������
$monitor($time,": ���� A:N1=%b N11=%b N24=%b N37=%b N50=%b N63=%b N76=%b N89=%b N102=%b    ���� B:N8=%b N21=%b N34=%b N47=%b N60=%b N73=%b N86=%b N99=%b N112=%b    ���� C:N14=%b N27=%b N40=%b N53=%b N66=%b N79=%b N92=%b N105=%b N115=%b    ���� E:N4=%b N17=%b N30=%b N43=%b N56=%b N69=%b N82=%b N95=%b N108=%b    �����:N223=%b N329=%b N370=%b N421=%b N430=%b N431=%b N432=%b",
tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115,tN4,tN17,tN30,tN43,tN56,tN69,tN82,tN95,tN108,tN223,tN329,tN370,tN421,tN430,tN431,tN432);

//�������� 1-�� ������������ � ��� ������������
#10;
     
     {tN1}=1'b0;
{tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN4}=1'b1;     
{tN17,tN30,tN43,tN56,tN69,tN82,tN95,tN108}=8'b00000000;      

//�������� 2-�� ������������ � ��� ������������
#10;
     
     {tN11}=1'b0;
{tN1,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN17}=1'b1;     
{tN4,tN30,tN43,tN56,tN69,tN82,tN95,tN108}=8'b00000000;

//�������� 3-�� ������������ � ��� ������������
#10;
     
     {tN24}=1'b0;
{tN1,tN11,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN30}=1'b1;     
{tN4,tN17,tN43,tN56,tN69,tN82,tN95,tN108}=8'b00000000;

//�������� 4-�� ������������ � ��� ������������
#10;
     
     {tN37}=1'b0;
{tN1,tN11,tN24,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN43}=1'b1;     
{tN4,tN17,tN30,tN56,tN69,tN82,tN95,tN108}=8'b00000000;

//�������� 5-�� ������������ � ��� ������������
#10;
     
     {tN50}=1'b0;
{tN1,tN11,tN24,tN37,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN56}=1'b1;     
{tN4,tN17,tN30,tN69,tN82,tN95,tN108}=8'b00000000;

//�������� 6-�� ������������ � ��� ������������
#10;
     
     {tN63}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN69}=1'b1;     
{tN4,tN17,tN30,tN43,tN56,tN82,tN95,tN108}=8'b00000000;


//�������� 7-�� ������������ � ��� ������������
#10;
     
     {tN76}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN82}=1'b1;     
{tN4,tN17,tN30,tN43,tN56,tN69,tN95,tN108}=8'b00000000;

//�������� 8-�� ������������ � ��� ������������
#10;
     
     {tN89}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN95}=1'b1;     
{tN4,tN17,tN30,tN43,tN56,tN69,tN82,tN108}=8'b00000000;

//�������� 9-�� ������������ � ��� ������������
#10;
     
     {tN102}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN108}=1'b1;     
{tN4,tN17,tN30,tN43,tN56,tN69,tN82,tN95}=8'b00000000;

//�������� 10-�� ������������ � ��� ������������
#10;
     
     {tN8}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN4}=1'b1;     
{tN17,tN30,tN43,tN56,tN69,tN82,tN95,tN108}=8'b00000000;      

//�������� 11-�� ������������ � ��� ������������
#10;
     
     {tN21}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN17}=1'b1;     
{tN4,tN30,tN43,tN56,tN69,tN82,tN95,tN108}=8'b00000000;

//�������� 12-�� ������������ � ��� ������������
#10;
     
     {tN34}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN30}=1'b1;     
{tN4,tN17,tN43,tN56,tN69,tN82,tN95,tN108}=8'b00000000;

//�������� 13-�� ������������ � ��� ������������
#10;
     
     {tN47}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN43}=1'b1;     
{tN4,tN17,tN30,tN56,tN69,tN82,tN95,tN108}=8'b00000000;

//�������� 14-�� ������������ � ��� ������������
#10;
     
     {tN60}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN56}=1'b1;     
{tN4,tN17,tN30,tN69,tN82,tN95,tN108}=8'b00000000;

//�������� 15-�� ������������ � ��� ������������
#10;
     
     {tN73}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN69}=1'b1;     
{tN4,tN17,tN30,tN43,tN56,tN82,tN95,tN108}=8'b00000000;


//�������� 16-�� ������������ � ��� ������������
#10;
     
     {tN86}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN82}=1'b1;     
{tN4,tN17,tN30,tN43,tN56,tN69,tN95,tN108}=8'b00000000;

//�������� 17-�� ������������ � ��� ������������
#10;
     
     {tN99}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN95}=1'b1;     
{tN4,tN17,tN30,tN43,tN56,tN69,tN82,tN108}=8'b00000000;

//�������� 18-�� ������������ � ��� ������������
#10;
     
     {tN112}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN108}=1'b1;     
{tN4,tN17,tN30,tN43,tN56,tN69,tN82,tN95}=8'b00000000;

//�������� 19-�� ������������ � ��� ������������
#10;
     
     {tN14}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN27,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN4}=1'b1;     
{tN17,tN30,tN43,tN56,tN69,tN82,tN95,tN108}=8'b00000000;      

//�������� 20-�� ������������ � ��� ������������
#10;
     
     {tN27}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN40,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN17}=1'b1;     
{tN4,tN30,tN43,tN56,tN69,tN82,tN95,tN108}=8'b00000000;

//�������� 21-�� ������������ � ��� ������������
#10;
     
     {tN40}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN53,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN30}=1'b1;     
{tN4,tN17,tN43,tN56,tN69,tN82,tN95,tN108}=8'b00000000;

//�������� 22-�� ������������ � ��� ������������
#10;
     
     {tN53}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN66,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN43}=1'b1;     
{tN4,tN17,tN30,tN56,tN69,tN82,tN95,tN108}=8'b00000000;

//�������� 23-�� ������������ � ��� ������������
#10;
     
     {tN66}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN79,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN56}=1'b1;     
{tN4,tN17,tN30,tN69,tN82,tN95,tN108}=8'b00000000;

//�������� 24-�� ������������ � ��� ������������
#10;
     
     {tN79}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN92,tN105,tN115}=26'b11111111111111111111111111;

     {tN69}=1'b1;     
{tN4,tN17,tN30,tN43,tN56,tN82,tN95,tN108}=8'b00000000;


//�������� 25-�� ������������ � ��� ������������
#10;
     
     {tN92}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN8,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN105,tN115}=26'b11111111111111111111111111;

     {tN82}=1'b1;     
{tN4,tN17,tN30,tN43,tN56,tN69,tN95,tN108}=8'b00000000;

//�������� 26-�� ������������ � ��� ������������
#10;
     
     {tN105}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN115}=26'b11111111111111111111111111;

     {tN95}=1'b1;     
{tN4,tN17,tN30,tN43,tN56,tN69,tN82,tN108}=8'b00000000;

//�������� 27-�� ������������ � ��� ������������
#10;
     
     {tN115}=1'b0;
{tN1,tN11,tN24,tN37,tN50,tN63,tN76,tN89,tN102,tN8,tN21,tN34,tN47,tN60,tN73,tN86,tN99,tN112,tN14,tN27,tN40,tN53,tN66,tN79,tN92,tN105}=26'b11111111111111111111111111;

     {tN108}=1'b1;     
{tN4,tN17,tN30,tN43,tN56,tN69,tN82,tN95}=8'b00000000;

end
endmodule