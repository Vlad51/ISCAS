
module c432 ( N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, 
        N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, 
        N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, 
        N421, N430, N431, N432 );
  input N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47,
         N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92,
         N95, N99, N102, N105, N108, N112, N115;
  output N223, N329, N370, N421, N430, N431, N432;
  wire   n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448;

  NAND2_X4 U185 ( .A1(N86), .A2(N329), .ZN(n184) );
  INV_X8 U186 ( .A(n184), .ZN(n265) );
  NOR2_X4 U187 ( .A1(N115), .A2(n439), .ZN(n185) );
  BUF_X8 U188 ( .A(n327), .Z(n186) );
  BUF_X8 U189 ( .A(N82), .Z(n187) );
  INV_X8 U190 ( .A(n264), .ZN(n188) );
  INV_X8 U191 ( .A(n188), .ZN(n189) );
  AND2_X4 U192 ( .A1(n336), .A2(n302), .ZN(n190) );
  AND2_X4 U193 ( .A1(n420), .A2(n270), .ZN(n191) );
  AND2_X4 U194 ( .A1(n256), .A2(n272), .ZN(n192) );
  NOR2_X4 U195 ( .A1(n194), .A2(n195), .ZN(n193) );
  INV_X8 U196 ( .A(n408), .ZN(n194) );
  INV_X8 U197 ( .A(n263), .ZN(n195) );
  BUF_X8 U198 ( .A(n345), .Z(n196) );
  BUF_X8 U199 ( .A(n331), .Z(n197) );
  NAND2_X4 U200 ( .A1(n322), .A2(n339), .ZN(n198) );
  NAND2_X4 U201 ( .A1(n336), .A2(n302), .ZN(n199) );
  BUF_X8 U202 ( .A(N63), .Z(n200) );
  BUF_X8 U203 ( .A(N69), .Z(n201) );
  NAND2_X4 U204 ( .A1(n366), .A2(n232), .ZN(n202) );
  BUF_X8 U205 ( .A(n330), .Z(n203) );
  BUF_X8 U206 ( .A(n322), .Z(n204) );
  NAND2_X4 U207 ( .A1(n199), .A2(n226), .ZN(n205) );
  BUF_X8 U208 ( .A(n340), .Z(n206) );
  INV_X8 U209 ( .A(n448), .ZN(n207) );
  INV_X8 U210 ( .A(n207), .ZN(n208) );
  BUF_X8 U211 ( .A(n344), .Z(n209) );
  BUF_X8 U212 ( .A(n342), .Z(n210) );
  NAND2_X4 U213 ( .A1(n355), .A2(n348), .ZN(n211) );
  NOR2_X4 U214 ( .A1(n198), .A2(n205), .ZN(n212) );
  NAND2_X4 U215 ( .A1(n425), .A2(n354), .ZN(n213) );
  NAND2_X4 U216 ( .A1(n295), .A2(n296), .ZN(n214) );
  INV_X8 U217 ( .A(n244), .ZN(n215) );
  NOR2_X4 U218 ( .A1(n317), .A2(n316), .ZN(n216) );
  NOR2_X4 U219 ( .A1(n350), .A2(n349), .ZN(n217) );
  OR2_X4 U220 ( .A1(n266), .A2(N14), .ZN(n218) );
  BUF_X8 U221 ( .A(n320), .Z(n219) );
  NOR2_X4 U222 ( .A1(n221), .A2(N102), .ZN(n220) );
  INV_X8 U223 ( .A(N108), .ZN(n221) );
  NAND2_X4 U224 ( .A1(n243), .A2(n241), .ZN(n222) );
  INV_X8 U225 ( .A(n222), .ZN(n296) );
  NAND2_X4 U226 ( .A1(n229), .A2(n210), .ZN(n223) );
  NAND2_X4 U227 ( .A1(n367), .A2(n279), .ZN(n224) );
  INV_X8 U228 ( .A(n224), .ZN(n325) );
  NAND2_X4 U229 ( .A1(n337), .A2(n226), .ZN(n225) );
  INV_X8 U230 ( .A(n259), .ZN(n226) );
  NAND2_X4 U231 ( .A1(n324), .A2(n325), .ZN(n227) );
  NAND2_X4 U232 ( .A1(n208), .A2(n203), .ZN(n228) );
  INV_X8 U233 ( .A(n207), .ZN(n229) );
  NOR2_X4 U234 ( .A1(n293), .A2(n292), .ZN(n230) );
  NAND2_X4 U235 ( .A1(n252), .A2(n217), .ZN(n231) );
  NOR2_X4 U236 ( .A1(n267), .A2(n218), .ZN(n232) );
  NAND2_X4 U237 ( .A1(n234), .A2(n263), .ZN(n233) );
  INV_X8 U238 ( .A(n233), .ZN(n245) );
  NOR2_X4 U239 ( .A1(n423), .A2(n422), .ZN(n234) );
  NAND2_X4 U240 ( .A1(n385), .A2(n386), .ZN(n235) );
  NAND2_X4 U241 ( .A1(n417), .A2(n392), .ZN(n236) );
  INV_X8 U242 ( .A(n236), .ZN(n264) );
  INV_X8 U243 ( .A(n247), .ZN(N329) );
  INV_X8 U244 ( .A(n247), .ZN(n238) );
  BUF_X8 U245 ( .A(N95), .Z(n239) );
  BUF_X8 U246 ( .A(N108), .Z(n240) );
  NAND2_X4 U247 ( .A1(n242), .A2(N69), .ZN(n241) );
  INV_X8 U248 ( .A(N63), .ZN(n242) );
  NAND2_X4 U249 ( .A1(n244), .A2(N82), .ZN(n243) );
  INV_X8 U250 ( .A(N76), .ZN(n244) );
  BUF_X8 U251 ( .A(n339), .Z(n246) );
  BUF_X8 U252 ( .A(n207), .Z(n247) );
  NAND2_X4 U253 ( .A1(n322), .A2(n339), .ZN(n248) );
  NAND2_X4 U254 ( .A1(n249), .A2(N82), .ZN(n327) );
  INV_X8 U255 ( .A(N86), .ZN(n249) );
  NOR2_X4 U256 ( .A1(n207), .A2(n190), .ZN(n250) );
  INV_X8 U257 ( .A(n250), .ZN(n370) );
  AND2_X4 U258 ( .A1(n326), .A2(n219), .ZN(n251) );
  NOR2_X4 U259 ( .A1(n335), .A2(n334), .ZN(n252) );
  NAND2_X4 U260 ( .A1(n230), .A2(n299), .ZN(n253) );
  NOR2_X4 U261 ( .A1(n248), .A2(n225), .ZN(n254) );
  NOR2_X4 U262 ( .A1(n264), .A2(n245), .ZN(n429) );
  NOR2_X4 U263 ( .A1(n255), .A2(N21), .ZN(n311) );
  INV_X8 U264 ( .A(n278), .ZN(n255) );
  INV_X8 U265 ( .A(N79), .ZN(n256) );
  NAND2_X4 U266 ( .A1(n257), .A2(n271), .ZN(n360) );
  INV_X8 U267 ( .A(N66), .ZN(n257) );
  NAND2_X4 U268 ( .A1(n187), .A2(n258), .ZN(n394) );
  NAND2_X4 U269 ( .A1(n215), .A2(n313), .ZN(n258) );
  NAND2_X4 U270 ( .A1(n260), .A2(n261), .ZN(n259) );
  NOR2_X4 U271 ( .A1(n305), .A2(n304), .ZN(n260) );
  NAND2_X4 U272 ( .A1(n309), .A2(n308), .ZN(n261) );
  AND2_X4 U273 ( .A1(n319), .A2(n327), .ZN(n307) );
  AND2_X4 U274 ( .A1(n262), .A2(n441), .ZN(n442) );
  OR2_X4 U275 ( .A1(n440), .A2(n439), .ZN(n262) );
  INV_X8 U276 ( .A(n424), .ZN(n263) );
  OR2_X4 U277 ( .A1(n266), .A2(n267), .ZN(n432) );
  INV_X8 U278 ( .A(N4), .ZN(n266) );
  AND2_X4 U279 ( .A1(N223), .A2(N1), .ZN(n267) );
  AND2_X4 U280 ( .A1(N43), .A2(n268), .ZN(n297) );
  INV_X8 U281 ( .A(N47), .ZN(n268) );
  AND2_X4 U282 ( .A1(N56), .A2(n269), .ZN(n310) );
  INV_X8 U283 ( .A(N60), .ZN(n269) );
  AND2_X4 U284 ( .A1(N43), .A2(n323), .ZN(n270) );
  AND2_X4 U285 ( .A1(N56), .A2(n321), .ZN(n271) );
  AND2_X4 U286 ( .A1(n343), .A2(n201), .ZN(n272) );
  AND2_X4 U287 ( .A1(n336), .A2(n239), .ZN(n273) );
  AND2_X4 U288 ( .A1(n272), .A2(n351), .ZN(n274) );
  INV_X8 U289 ( .A(n431), .ZN(N370) );
  BUF_X8 U290 ( .A(N30), .Z(n276) );
  BUF_X8 U291 ( .A(N11), .Z(n277) );
  BUF_X8 U292 ( .A(N17), .Z(n278) );
  NAND2_X4 U293 ( .A1(n359), .A2(n280), .ZN(n279) );
  INV_X8 U294 ( .A(n360), .ZN(n280) );
  INV_X8 U295 ( .A(N30), .ZN(n281) );
  NOR2_X4 U296 ( .A1(n281), .A2(N24), .ZN(n284) );
  INV_X8 U297 ( .A(N17), .ZN(n282) );
  NOR2_X4 U298 ( .A1(n282), .A2(N11), .ZN(n283) );
  NOR2_X4 U299 ( .A1(n284), .A2(n283), .ZN(n287) );
  INV_X8 U300 ( .A(N1), .ZN(n285) );
  NAND2_X4 U301 ( .A1(N4), .A2(n285), .ZN(n286) );
  NAND2_X4 U302 ( .A1(n287), .A2(n286), .ZN(n293) );
  INV_X8 U303 ( .A(N37), .ZN(n288) );
  NAND2_X4 U304 ( .A1(N43), .A2(n288), .ZN(n291) );
  INV_X8 U305 ( .A(N50), .ZN(n289) );
  NAND2_X4 U306 ( .A1(N56), .A2(n289), .ZN(n290) );
  NAND2_X4 U307 ( .A1(n291), .A2(n290), .ZN(n292) );
  NOR2_X4 U308 ( .A1(n293), .A2(n292), .ZN(n309) );
  INV_X8 U309 ( .A(n201), .ZN(n312) );
  INV_X8 U310 ( .A(n240), .ZN(n298) );
  INV_X8 U311 ( .A(N95), .ZN(n301) );
  NOR2_X4 U312 ( .A1(n301), .A2(N89), .ZN(n294) );
  NOR2_X4 U313 ( .A1(n294), .A2(n220), .ZN(n295) );
  NAND2_X4 U314 ( .A1(n296), .A2(n295), .ZN(n306) );
  INV_X8 U315 ( .A(n306), .ZN(n299) );
  NAND2_X4 U316 ( .A1(n230), .A2(n299), .ZN(N223) );
  NAND2_X4 U317 ( .A1(n313), .A2(N37), .ZN(n323) );
  NAND2_X4 U318 ( .A1(n323), .A2(n297), .ZN(n322) );
  NOR2_X4 U319 ( .A1(n298), .A2(N112), .ZN(n300) );
  NAND2_X4 U320 ( .A1(n299), .A2(n309), .ZN(n313) );
  NAND2_X4 U321 ( .A1(n253), .A2(N102), .ZN(n340) );
  NAND2_X4 U322 ( .A1(n340), .A2(n300), .ZN(n339) );
  NOR2_X4 U323 ( .A1(n301), .A2(N99), .ZN(n302) );
  NAND2_X4 U324 ( .A1(N223), .A2(N89), .ZN(n336) );
  NAND2_X4 U325 ( .A1(n336), .A2(n302), .ZN(n337) );
  INV_X8 U326 ( .A(N8), .ZN(n303) );
  NAND2_X4 U327 ( .A1(n303), .A2(N4), .ZN(n319) );
  NOR2_X4 U328 ( .A1(n319), .A2(N1), .ZN(n305) );
  NOR2_X4 U329 ( .A1(n327), .A2(n215), .ZN(n304) );
  NOR2_X4 U330 ( .A1(n307), .A2(n214), .ZN(n308) );
  NAND2_X4 U331 ( .A1(n253), .A2(N50), .ZN(n321) );
  NAND2_X4 U332 ( .A1(n310), .A2(n321), .ZN(n320) );
  NAND2_X4 U333 ( .A1(n313), .A2(n277), .ZN(n331) );
  NAND2_X4 U334 ( .A1(n331), .A2(n311), .ZN(n330) );
  NAND2_X4 U335 ( .A1(n320), .A2(n330), .ZN(n317) );
  NOR2_X4 U336 ( .A1(n312), .A2(N73), .ZN(n314) );
  NAND2_X4 U337 ( .A1(n253), .A2(n200), .ZN(n343) );
  NAND2_X4 U338 ( .A1(n343), .A2(n314), .ZN(n342) );
  NOR2_X4 U339 ( .A1(n281), .A2(N34), .ZN(n315) );
  NAND2_X4 U340 ( .A1(N223), .A2(N24), .ZN(n345) );
  NAND2_X4 U341 ( .A1(n345), .A2(n315), .ZN(n344) );
  NAND2_X4 U342 ( .A1(n342), .A2(n344), .ZN(n316) );
  NOR2_X4 U343 ( .A1(n317), .A2(n316), .ZN(n318) );
  NAND2_X4 U344 ( .A1(n318), .A2(n254), .ZN(n448) );
  NAND2_X4 U345 ( .A1(n216), .A2(n212), .ZN(n326) );
  NAND2_X4 U346 ( .A1(n326), .A2(n319), .ZN(n366) );
  INV_X8 U347 ( .A(N14), .ZN(n430) );
  NAND2_X4 U348 ( .A1(n326), .A2(n219), .ZN(n359) );
  NAND2_X4 U349 ( .A1(n208), .A2(n204), .ZN(n377) );
  INV_X8 U350 ( .A(N53), .ZN(n420) );
  NAND2_X4 U351 ( .A1(n377), .A2(n191), .ZN(n324) );
  NAND2_X4 U352 ( .A1(n325), .A2(n324), .ZN(n335) );
  NOR2_X4 U353 ( .A1(n394), .A2(N92), .ZN(n329) );
  NAND2_X4 U354 ( .A1(n326), .A2(n186), .ZN(n328) );
  NAND2_X4 U355 ( .A1(n329), .A2(n328), .ZN(n356) );
  NAND2_X4 U356 ( .A1(n197), .A2(n278), .ZN(n388) );
  NOR2_X4 U357 ( .A1(n388), .A2(N27), .ZN(n332) );
  NAND2_X4 U358 ( .A1(n228), .A2(n332), .ZN(n333) );
  NAND2_X4 U359 ( .A1(n356), .A2(n333), .ZN(n334) );
  NOR2_X4 U360 ( .A1(n227), .A2(n334), .ZN(n419) );
  INV_X8 U361 ( .A(N105), .ZN(n396) );
  NAND2_X4 U362 ( .A1(n396), .A2(n273), .ZN(n371) );
  INV_X8 U363 ( .A(n371), .ZN(n338) );
  NAND2_X4 U364 ( .A1(n370), .A2(n338), .ZN(n341) );
  NAND2_X4 U365 ( .A1(n229), .A2(n246), .ZN(n364) );
  NAND2_X4 U366 ( .A1(n206), .A2(n240), .ZN(n439) );
  NAND2_X4 U367 ( .A1(n365), .A2(n341), .ZN(n350) );
  NAND2_X4 U368 ( .A1(n229), .A2(n209), .ZN(n347) );
  NAND2_X4 U369 ( .A1(n196), .A2(n276), .ZN(n380) );
  NOR2_X4 U370 ( .A1(n380), .A2(N40), .ZN(n346) );
  NAND2_X4 U371 ( .A1(n347), .A2(n346), .ZN(n348) );
  NAND2_X4 U372 ( .A1(n355), .A2(n348), .ZN(n349) );
  NOR2_X4 U373 ( .A1(n350), .A2(n211), .ZN(n421) );
  NAND2_X4 U374 ( .A1(N73), .A2(N329), .ZN(n351) );
  NAND2_X4 U375 ( .A1(N370), .A2(N79), .ZN(n352) );
  NAND2_X4 U376 ( .A1(n352), .A2(n274), .ZN(n412) );
  NAND2_X4 U377 ( .A1(N60), .A2(N329), .ZN(n353) );
  NAND2_X4 U378 ( .A1(n271), .A2(n353), .ZN(n426) );
  INV_X8 U379 ( .A(n426), .ZN(n354) );
  NAND2_X4 U380 ( .A1(n252), .A2(n421), .ZN(n391) );
  NAND2_X4 U381 ( .A1(n391), .A2(N66), .ZN(n425) );
  NAND2_X4 U382 ( .A1(n425), .A2(n354), .ZN(n409) );
  NAND2_X4 U383 ( .A1(n223), .A2(n192), .ZN(n355) );
  INV_X8 U384 ( .A(N40), .ZN(n378) );
  NOR2_X4 U385 ( .A1(n355), .A2(n378), .ZN(n358) );
  NOR2_X4 U386 ( .A1(n356), .A2(n378), .ZN(n357) );
  NOR2_X4 U387 ( .A1(n358), .A2(n357), .ZN(n363) );
  NOR2_X4 U388 ( .A1(n251), .A2(n360), .ZN(n361) );
  NAND2_X4 U389 ( .A1(N40), .A2(n361), .ZN(n362) );
  NAND2_X4 U390 ( .A1(n363), .A2(n362), .ZN(n376) );
  NAND2_X4 U391 ( .A1(n364), .A2(n185), .ZN(n365) );
  NOR2_X4 U392 ( .A1(n365), .A2(n378), .ZN(n369) );
  NAND2_X4 U393 ( .A1(n366), .A2(n232), .ZN(n367) );
  NOR2_X4 U394 ( .A1(n202), .A2(n378), .ZN(n368) );
  NOR2_X4 U395 ( .A1(n369), .A2(n368), .ZN(n374) );
  NOR2_X4 U396 ( .A1(n250), .A2(n371), .ZN(n372) );
  NAND2_X4 U397 ( .A1(N40), .A2(n372), .ZN(n373) );
  NAND2_X4 U398 ( .A1(n374), .A2(n373), .ZN(n375) );
  NOR2_X4 U399 ( .A1(n376), .A2(n375), .ZN(n386) );
  NAND2_X4 U400 ( .A1(n377), .A2(n191), .ZN(n379) );
  NOR2_X4 U401 ( .A1(n379), .A2(n378), .ZN(n384) );
  INV_X8 U402 ( .A(n380), .ZN(n382) );
  NAND2_X4 U403 ( .A1(N34), .A2(n238), .ZN(n381) );
  NAND2_X4 U404 ( .A1(n382), .A2(n381), .ZN(n383) );
  NOR2_X4 U405 ( .A1(n384), .A2(n383), .ZN(n385) );
  NAND2_X4 U406 ( .A1(n385), .A2(n386), .ZN(n401) );
  NAND2_X4 U407 ( .A1(n213), .A2(n235), .ZN(n387) );
  NOR2_X4 U408 ( .A1(n412), .A2(n387), .ZN(n393) );
  INV_X8 U409 ( .A(n388), .ZN(n390) );
  NAND2_X4 U410 ( .A1(N21), .A2(N329), .ZN(n389) );
  NAND2_X4 U411 ( .A1(n390), .A2(n389), .ZN(n418) );
  INV_X8 U412 ( .A(n418), .ZN(n392) );
  NAND2_X4 U413 ( .A1(n231), .A2(N27), .ZN(n417) );
  NOR2_X4 U414 ( .A1(n393), .A2(n189), .ZN(n407) );
  INV_X8 U415 ( .A(n401), .ZN(n427) );
  NOR2_X4 U416 ( .A1(n265), .A2(n394), .ZN(n436) );
  NAND2_X4 U417 ( .A1(n231), .A2(N92), .ZN(n395) );
  NAND2_X4 U418 ( .A1(n395), .A2(n436), .ZN(n411) );
  INV_X8 U419 ( .A(n391), .ZN(n431) );
  NOR2_X4 U420 ( .A1(n431), .A2(n396), .ZN(n398) );
  NAND2_X4 U421 ( .A1(N99), .A2(N329), .ZN(n397) );
  NAND2_X4 U422 ( .A1(n273), .A2(n397), .ZN(n441) );
  NOR2_X4 U423 ( .A1(n398), .A2(n441), .ZN(n399) );
  NAND2_X4 U424 ( .A1(n399), .A2(n411), .ZN(n400) );
  NOR2_X4 U425 ( .A1(n400), .A2(n427), .ZN(n405) );
  NAND2_X4 U426 ( .A1(n231), .A2(N53), .ZN(n408) );
  NAND2_X4 U427 ( .A1(n235), .A2(n408), .ZN(n403) );
  NAND2_X4 U428 ( .A1(N47), .A2(n238), .ZN(n402) );
  NAND2_X4 U429 ( .A1(n270), .A2(n402), .ZN(n424) );
  NOR2_X4 U430 ( .A1(n403), .A2(n424), .ZN(n404) );
  NOR2_X4 U431 ( .A1(n405), .A2(n404), .ZN(n406) );
  NAND2_X4 U432 ( .A1(n406), .A2(n407), .ZN(N432) );
  INV_X8 U433 ( .A(n409), .ZN(n410) );
  NOR2_X4 U434 ( .A1(n193), .A2(n410), .ZN(n414) );
  NAND2_X4 U435 ( .A1(n412), .A2(n411), .ZN(n413) );
  NAND2_X4 U436 ( .A1(n414), .A2(n413), .ZN(n416) );
  NOR2_X4 U437 ( .A1(n189), .A2(n427), .ZN(n415) );
  NAND2_X4 U438 ( .A1(n416), .A2(n415), .ZN(N431) );
  NOR2_X4 U439 ( .A1(n419), .A2(n420), .ZN(n423) );
  NOR2_X4 U440 ( .A1(n217), .A2(n420), .ZN(n422) );
  NOR2_X4 U441 ( .A1(n410), .A2(n427), .ZN(n428) );
  NAND2_X4 U442 ( .A1(n429), .A2(n428), .ZN(N430) );
  NOR2_X4 U443 ( .A1(n431), .A2(n430), .ZN(n433) );
  NOR2_X4 U444 ( .A1(n433), .A2(n432), .ZN(n435) );
  NAND2_X4 U445 ( .A1(N8), .A2(N329), .ZN(n434) );
  NAND2_X4 U446 ( .A1(n435), .A2(n434), .ZN(n445) );
  NAND2_X4 U447 ( .A1(N430), .A2(n445), .ZN(n447) );
  NOR2_X4 U448 ( .A1(n436), .A2(n274), .ZN(n443) );
  INV_X8 U449 ( .A(n238), .ZN(n438) );
  INV_X8 U450 ( .A(N112), .ZN(n437) );
  NOR2_X4 U451 ( .A1(n438), .A2(n437), .ZN(n440) );
  NAND2_X4 U452 ( .A1(n443), .A2(n442), .ZN(n444) );
  NAND2_X4 U453 ( .A1(n444), .A2(n445), .ZN(n446) );
  NAND2_X4 U454 ( .A1(n447), .A2(n446), .ZN(N421) );
endmodule

