//  file :c432.v
// Verilog 
// c432 
// Ninputs 36 
// Noutputs 7 
// NtotalGates 160 
// NOT1 40 
// NAND2 64 
// NOR2 19 
// AND9 3 
// XOR2 18 
// NAND4 14 
// AND8 1 
// NAND3 1 
 
module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30, 
N34,N37,N40,N43,N47,N50,N53,N56,N60,N63, 
N66,N69,N73,N76,N79,N82,N86,N89,N92,N95, 
N99,N102,N105,N108,N112,N115,N223,N329,N370,N421, 
N430,N431,N432); 
 
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30, 
N34,N37,N40,N43,N47,N50,N53,N56,N60,N63, 
N66,N69,N73,N76,N79,N82,N86,N89,N92,N95, 
N99,N102,N105,N108,N112,N115; 
 
output N223,N329,N370,N421,N430,N431,N432; 
 
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135, 
N138,N139,N142,N143,N146,N147,N150,N151,N154,N157, 
N158,N159,N162,N165,N168,N171,N174,N177,N180,N183, 
N184,N185,N186,N187,N188,N189,N190,N191,N192,N193, 
N194,N195,N196,N197,N198,N199,N203,N213,N224,N227, 
N230,N233,N236,N239,N242,N243,N246,N247,N250,N251, 
N254,N255,N256,N257,N258,N259,N260,N263,N264,N267, 
N270,N273,N276,N279,N282,N285,N288,N289,N290,N291, 
N292,N293,N294,N295,N296,N300,N301,N302,N303,N304, 
N305,N306,N307,N308,N309,N319,N330,N331,N332,N333, 
N334,N335,N336,N337,N338,N339,N340,N341,N342,N343, 
N344,N345,N346,N347,N348,N349,N350,N351,N352,N353, 
N354,N355,N356,N357,N360,N371,N372,N373,N374,N375, 
N376,N377,N378,N379,N380,N381,N386,N393,N399,N404, 
N407,N411,N414,N415,N416,N417,N418,N419,N420,N422, 
N425,N428,N429; 
  IN1 NOT1_1  (  .Q(N118), .A(N1) ); 
  IN1 NOT1_2  (  .Q(N119), .A(N4) ); 
  IN1 NOT1_3  (  .Q(N122), .A(N11) ); 
  IN1 NOT1_4  (  .Q(N123), .A(N17) ); 
  IN1 NOT1_5  (  .Q(N126), .A(N24) ); 
  IN1 NOT1_6  (  .Q(N127), .A(N30) ); 
  IN1 NOT1_7  (  .Q(N130), .A(N37) ); 
  IN1 NOT1_8  (  .Q(N131), .A(N43) ); 
  IN1 NOT1_9  (  .Q(N134), .A(N50) ); 
  IN1 NOT1_10  (  .Q(N135), .A(N56) ); 
  IN1 NOT1_11  (  .Q(N138), .A(N63) ); 
  IN1 NOT1_12  (  .Q(N139), .A(N69) ); 
  IN1 NOT1_13  (  .Q(N142), .A(N76) ); 
  IN1 NOT1_14  (  .Q(N143), .A(N82) ); 
  IN1 NOT1_15  (  .Q(N146), .A(N89) ); 
  IN1 NOT1_16  (  .Q(N147), .A(N95) ); 
  IN1 NOT1_17  (  .Q(N150), .A(N102) ); 
  IN1 NOT1_18  (  .Q(N151), .A(N108) ); 
  NA2 NAND2_19  (  .Q(N154), .A(N118), .B(N4) ); 
  NO2 NOR2_20  (  .Q(N157), .A(N8), .B(N119) ); 
  NO2 NOR2_21  (  .Q(N158), .A(N14), .B(N119) ); 
  NA2 NAND2_22  (  .Q(N159), .A(N122), .B(N17) ); 
  NA2 NAND2_23  (  .Q(N162), .A(N126), .B(N30) ); 
  NA2 NAND2_24  (  .Q(N165), .A(N130), .B(N43) ); 
  NA2 NAND2_25  (  .Q(N168), .A(N134), .B(N56) ); 
  NA2 NAND2_26  (  .Q(N171), .A(N138), .B(N69) ); 
  NA2 NAND2_27  (  .Q(N174), .A(N142), .B(N82) ); 
  NA2 NAND2_28  (  .Q(N177), .A(N146), .B(N95) ); 
  NA2 NAND2_29  (  .Q(N180), .A(N150), .B(N108) ); 
  NO2 NOR2_30  (  .Q(N183), .A(N21), .B(N123) ); 
  NO2 NOR2_31  (  .Q(N184), .A(N27), .B(N123) ); 
  NO2 NOR2_32  (  .Q(N185), .A(N34), .B(N127) ); 
  NO2 NOR2_33  (  .Q(N186), .A(N40), .B(N127) ); 
  NO2 NOR2_34  (  .Q(N187), .A(N47), .B(N131) ); 
  NO2 NOR2_35  (  .Q(N188), .A(N53), .B(N131) ); 
  NO2 NOR2_36  (  .Q(N189), .A(N60), .B(N135) ); 
  NO2 NOR2_37  (  .Q(N190), .A(N66), .B(N135) ); 
  NO2 NOR2_38  (  .Q(N191), .A(N73), .B(N139) ); 
  NO2 NOR2_39  (  .Q(N192), .A(N79), .B(N139) ); 
  NO2 NOR2_40  (  .Q(N193), .A(N86), .B(N143) ); 
  NO2 NOR2_41  (  .Q(N194), .A(N92), .B(N143) ); 
  NO2 NOR2_42  (  .Q(N195), .A(N99), .B(N147) ); 
  NO2 NOR2_43  (  .Q(N196), .A(N105), .B(N147) ); 
  NO2 NOR2_44  (  .Q(N197), .A(N112), .B(N151) ); 
  NO2 NOR2_45  (  .Q(N198), .A(N115), .B(N151) ); 
  AND9 AND9_46  (  .Q(N199), .A(N154), .B(N159), .C(N162), .D(N165), .E(N168), .F(N171), .G(N174), .H(N177), .I(N180) ); 
  IN1 NOT1_47  (  .Q(N203), .A(N199) ); 
  IN1 NOT1_48  (  .Q(N213), .A(N199) ); 
  IN1 NOT1_49  (  .Q(N223), .A(N199) ); 
  EO1 XOR2_50  (  .Q(N224), .A(N203), .B(N154) ); 
  EO1 XOR2_51  (  .Q(N227), .A(N203), .B(N159) ); 
  EO1 XOR2_52  (  .Q(N230), .A(N203), .B(N162) ); 
  EO1 XOR2_53  (  .Q(N233), .A(N203), .B(N165) ); 
  EO1 XOR2_54  (  .Q(N236), .A(N203), .B(N168) ); 
  EO1 XOR2_55  (  .Q(N239), .A(N203), .B(N171) ); 
  NA2 NAND2_56  (  .Q(N242), .A(N1), .B(N213) ); 
  EO1 XOR2_57  (  .Q(N243), .A(N203), .B(N174) ); 
  NA2 NAND2_58  (  .Q(N246), .A(N213), .B(N11) ); 
  EO1 XOR2_59  (  .Q(N247), .A(N203), .B(N177) ); 
  NA2 NAND2_60  (  .Q(N250), .A(N213), .B(N24) ); 
  EO1 XOR2_61  (  .Q(N251), .A(N203), .B(N180) ); 
  NA2 NAND2_62  (  .Q(N254), .A(N213), .B(N37) ); 
  NA2 NAND2_63  (  .Q(N255), .A(N213), .B(N50) ); 
  NA2 NAND2_64  (  .Q(N256), .A(N213), .B(N63) ); 
  NA2 NAND2_65  (  .Q(N257), .A(N213), .B(N76) ); 
  NA2 NAND2_66  (  .Q(N258), .A(N213), .B(N89) ); 
  NA2 NAND2_67  (  .Q(N259), .A(N213), .B(N102) ); 
  NA2 NAND2_68  (  .Q(N260), .A(N224), .B(N157) ); 
  NA2 NAND2_69  (  .Q(N263), .A(N224), .B(N158) ); 
  NA2 NAND2_70  (  .Q(N264), .A(N227), .B(N183) ); 
  NA2 NAND2_71  (  .Q(N267), .A(N230), .B(N185) ); 
  NA2 NAND2_72  (  .Q(N270), .A(N233), .B(N187) ); 
  NA2 NAND2_73  (  .Q(N273), .A(N236), .B(N189) ); 
  NA2 NAND2_74  (  .Q(N276), .A(N239), .B(N191) ); 
  NA2 NAND2_75  (  .Q(N279), .A(N243), .B(N193) ); 
  NA2 NAND2_76  (  .Q(N282), .A(N247), .B(N195) ); 
  NA2 NAND2_77  (  .Q(N285), .A(N251), .B(N197) ); 
  NA2 NAND2_78  (  .Q(N288), .A(N227), .B(N184) ); 
  NA2 NAND2_79  (  .Q(N289), .A(N230), .B(N186) ); 
  NA2 NAND2_80  (  .Q(N290), .A(N233), .B(N188) ); 
  NA2 NAND2_81  (  .Q(N291), .A(N236), .B(N190) ); 
  NA2 NAND2_82  (  .Q(N292), .A(N239), .B(N192) ); 
  NA2 NAND2_83  (  .Q(N293), .A(N243), .B(N194) ); 
  NA2 NAND2_84  (  .Q(N294), .A(N247), .B(N196) ); 
  NA2 NAND2_85  (  .Q(N295), .A(N251), .B(N198) ); 
  AND9 AND9_86  (  .Q(N296), .A(N260), .B(N264), .C(N267), .D(N270), .E(N273), .F(N276), .G(N279), .H(N282), .I(N285) ); 
  IN1 NOT1_87  (  .Q(N300), .A(N263) ); 
  IN1 NOT1_88  (  .Q(N301), .A(N288) ); 
  IN1 NOT1_89  (  .Q(N302), .A(N289) ); 
  IN1 NOT1_90  (  .Q(N303), .A(N290) ); 
  IN1 NOT1_91  (  .Q(N304), .A(N291) ); 
  IN1 NOT1_92  (  .Q(N305), .A(N292) ); 
  IN1 NOT1_93  (  .Q(N306), .A(N293) ); 
  IN1 NOT1_94  (  .Q(N307), .A(N294) ); 
  IN1 NOT1_95  (  .Q(N308), .A(N295) ); 
  IN1 NOT1_96  (  .Q(N309), .A(N296) ); 
  IN1 NOT1_97  (  .Q(N319), .A(N296) ); 
  IN1 NOT1_98  (  .Q(N329), .A(N296) ); 
  EO1 XOR2_99  (  .Q(N330), .A(N309), .B(N260) ); 
  EO1 XOR2_100  (  .Q(N331), .A(N309), .B(N264) ); 
  EO1 XOR2_101  (  .Q(N332), .A(N309), .B(N267) ); 
  EO1 XOR2_102  (  .Q(N333), .A(N309), .B(N270) ); 
  NA2 NAND2_103  (  .Q(N334), .A(N8), .B(N319) ); 
  EO1 XOR2_104  (  .Q(N335), .A(N309), .B(N273) ); 
  NA2 NAND2_105  (  .Q(N336), .A(N319), .B(N21) ); 
  EO1 XOR2_106  (  .Q(N337), .A(N309), .B(N276) ); 
  NA2 NAND2_107  (  .Q(N338), .A(N319), .B(N34) ); 
  EO1 XOR2_108  (  .Q(N339), .A(N309), .B(N279) ); 
  NA2 NAND2_109  (  .Q(N340), .A(N319), .B(N47) ); 
  EO1 XOR2_110  (  .Q(N341), .A(N309), .B(N282) ); 
  NA2 NAND2_111  (  .Q(N342), .A(N319), .B(N60) ); 
  EO1 XOR2_112  (  .Q(N343), .A(N309), .B(N285) ); 
  NA2 NAND2_113  (  .Q(N344), .A(N319), .B(N73) ); 
  NA2 NAND2_114  (  .Q(N345), .A(N319), .B(N86) ); 
  NA2 NAND2_115  (  .Q(N346), .A(N319), .B(N99) ); 
  NA2 NAND2_116  (  .Q(N347), .A(N319), .B(N112) ); 
  NA2 NAND2_117  (  .Q(N348), .A(N330), .B(N300) ); 
  NA2 NAND2_118  (  .Q(N349), .A(N331), .B(N301) ); 
  NA2 NAND2_119  (  .Q(N350), .A(N332), .B(N302) ); 
  NA2 NAND2_120  (  .Q(N351), .A(N333), .B(N303) ); 
  NA2 NAND2_121  (  .Q(N352), .A(N335), .B(N304) ); 
  NA2 NAND2_122  (  .Q(N353), .A(N337), .B(N305) ); 
  NA2 NAND2_123  (  .Q(N354), .A(N339), .B(N306) ); 
  NA2 NAND2_124  (  .Q(N355), .A(N341), .B(N307) ); 
  NA2 NAND2_125  (  .Q(N356), .A(N343), .B(N308) ); 
  AND9 AND9_126  (  .Q(N357), .A(N348), .B(N349), .C(N350), .D(N351), .E(N352), .F(N353), .G(N354), .H(N355), .I(N356) ); 
  IN1 NOT1_127  (  .Q(N360), .A(N357) ); 
  IN1 NOT1_128  (  .Q(N370), .A(N357) ); 
  NA2 NAND2_129  (  .Q(N371), .A(N14), .B(N360) ); 
  NA2 NAND2_130  (  .Q(N372), .A(N360), .B(N27) ); 
  NA2 NAND2_131  (  .Q(N373), .A(N360), .B(N40) ); 
  NA2 NAND2_132  (  .Q(N374), .A(N360), .B(N53) ); 
  NA2 NAND2_133  (  .Q(N375), .A(N360), .B(N66) ); 
  NA2 NAND2_134  (  .Q(N376), .A(N360), .B(N79) ); 
  NA2 NAND2_135  (  .Q(N377), .A(N360), .B(N92) ); 
  NA2 NAND2_136  (  .Q(N378), .A(N360), .B(N105) ); 
  NA2 NAND2_137  (  .Q(N379), .A(N360), .B(N115) ); 
  NA4 NAND4_138  (  .Q(N380), .A(N4), .B(N242), .C(N334), .D(N371) ); 
  NA4 NAND4_139  (  .Q(N381), .A(N246), .B(N336), .C(N372), .D(N17) ); 
  NA4 NAND4_140  (  .Q(N386), .A(N250), .B(N338), .C(N373), .D(N30) ); 
  NA4 NAND4_141  (  .Q(N393), .A(N254), .B(N340), .C(N374), .D(N43) ); 
  NA4 NAND4_142  (  .Q(N399), .A(N255), .B(N342), .C(N375), .D(N56) ); 
  NA4 NAND4_143  (  .Q(N404), .A(N256), .B(N344), .C(N376), .D(N69) ); 
  NA4 NAND4_144  (  .Q(N407), .A(N257), .B(N345), .C(N377), .D(N82) ); 
  NA4 NAND4_145  (  .Q(N411), .A(N258), .B(N346), .C(N378), .D(N95) ); 
  NA4 NAND4_146  (  .Q(N414), .A(N259), .B(N347), .C(N379), .D(N108) ); 
  IN1 NOT1_147  (  .Q(N415), .A(N380) ); 
  AND8 AND8_148  (  .Q(N416), .A(N381), .B(N386), .C(N393), .D(N399), .E(N404), .F(N407), .G(N411), .H(N414) ); 
  IN1 NOT1_149  (  .Q(N417), .A(N393) ); 
  IN1 NOT1_150  (  .Q(N418), .A(N404) ); 
  IN1 NOT1_151  (  .Q(N419), .A(N407) ); 
  IN1 NOT1_152  (  .Q(N420), .A(N411) ); 
  NO2 NOR2_153  (  .Q(N421), .A(N415), .B(N416) ); 
  NA2 NAND2_154  (  .Q(N422), .A(N386), .B(N417) ); 
  NA4 NAND4_155  (  .Q(N425), .A(N386), .B(N393), .C(N418), .D(N399) ); 
  NA3 NAND3_156  (  .Q(N428), .A(N399), .B(N393), .C(N419) ); 
  NA4 NAND4_157  (  .Q(N429), .A(N386), .B(N393), .C(N407), .D(N420) ); 
  NA4 NAND4_158  (  .Q(N430), .A(N381), .B(N386), .C(N422), .D(N399) ); 
  NA4 NAND4_159  (  .Q(N431), .A(N381), .B(N386), .C(N425), .D(N428) ); 
  NA4 NAND4_160  (  .Q(N432), .A(N381), .B(N422), .C(N425), .D(N429) ); 
endmodule 
