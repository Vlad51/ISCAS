HEADER $
    CIRCUIT NAME $
         c17 $                     
    TECHNOLOGY $
         ECL $
    LAST UPDATE $
         Jan 21, 1985 $

PARTS $
    A6     NAND/2 $
    A7     NAND/2 $
    A8     NAND/2 $
    A9     NAND/2 $
    A10    NAND/2 $
    A11    NAND/2 $

CONNECTIONS $
         A1       A6.1     $
         A3       A6.2     A7.1     $
         A6       A6.3     A10.1    $
         A4       A7.2     $
         A7       A7.3     A8.2     A9.1     $
         A2       A8.1     $
         A8       A8.3     A10.2    A11.1    $
         A5       A9.2     $
         A9       A9.3     A11.2    $
         A10      A10.3    $
         A11      A11.3    $

EXTERNALS $
         A1       $
         A2       $
         A3       $
         A4       $
         A5       $
         A10      $
         A11      $

END $
